module or_gate(out, a, b);
input a, b;
output out;
or(out, a, b);
endmodule
